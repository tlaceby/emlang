module compiler

import frontend.parser.lexer { SourceFile }
import frontend.parser { Parser }
import vm.values { CodeVal }
import time
import frontend.analysis


// EMCompiler is responsible for taking an abstract syntax tree (AST) and generating
// bytecode for the given program.
pub struct EMCompiler {
	mut:
	parser Parser     // The parser to produce the AST from the source code
	code CodeVal      // The generated bytecode
}

// emit_bytecode takes a source file and produces the bytecode for it.
pub fn (mut c EMCompiler) emit_bytecode (entry SourceFile) CodeVal {
	start := time.now()
	ast := c.parser.produce_ast(entry)
	mut checker := analysis.TypeChecker{}
	checker.perform_type_analysis(ast)
	// println(ast)
	end := time.now()

	println("time: ${end - start}")
	return c.code
}
